module xor_gate_1bit(
	output result,
	input A,
	input B
);
	xor xor_gate(result, A, B);
	
endmodule

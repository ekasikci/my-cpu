module or_gate_1bit(
	output result,
	input A,
	input B
);
	or or_gate(result, A, B);
	
endmodule
